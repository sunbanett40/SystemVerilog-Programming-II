    Mac OS X            	   2  d     �                                      ATTR      �     �                      com.apple.TextEncoding          com.apple.lastuseddate#PS      '   S  com.dropbox.attributes     z     com.dropbox.attrs    UTF-8;134217984F=�[    +��     x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK��4�bG#� #?ǲ$w�rC�2�t[[���Z ���

��Y�%\      ���ゅ